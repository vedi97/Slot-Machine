/******************************************************************
***Desiged by:		Vedi Ghahremanyans			                      ***
***Topic:		ECE 526 Final Project			                          ***
***Project Name:	Basic Slot Machine			                      ***
***								                                              ***
***File Name: 		rgen1.v					                              ***
*******************************************************************
***rgen1 module will take the seed1 generated by the hardware	  ***			
***and put in the random1 register in order to do logical	      ***
***operation to create random #1.				                        ***
*******************************************************************/		
`timescale 1 ns / 1 ns

module rgen1(clk, rnum1, seed1);

//**************INPUT/OUTPUT**************
	input  clk;
	input  [5:0] seed1;
	output [3:0] rnum1;
//**************INPUT/OUTPUT**************



//**************Register**************
	reg [5:0] random1;
//**************Register**************



//**************Functionality**************
	always @(posedge clk)
		begin
			random1 = seed1;
			random1[0] <= random1[4] ^ random1[5];
			random1[5:1] <= random1[4:0];
		end

	assign rnum1 = random1[3:0];
//**************Functionality**************

endmodule
