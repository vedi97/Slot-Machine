/******************************************************************
***Desiged by:		Vedi Ghahremanyans			***
***Topic:		ECE 526 Final Project			***
***Project Name:	Basic Slot Machine			***
***								***
***File Name: 		RandomNumberHandler.v			***
*******************************************************************
***RandomNumberHandler will generate rnum1, rnum2, and rnum3 by ***			
***using seed1, seed2, and seed3 generated by the hardware 	***
***and decided if $1 or $2 wins or not. 			***
*******************************************************************/		
`timescale 1 ns / 1 ns

module RandomNumberHandler(clk, rnum1, rnum2, rnum3, seed1, seed2, seed3, bet_1d, bet_2d);


//**************Parameters**************
parameter [1:0]one_d_win	= 2'b00;	//Binary Code to win if $1 is bet
parameter [1:0]one_d_lose	= 2'b01;	//Binary Code to lose  if $1 is bet
parameter [1:0]two_d_win 	= 2'b10;	//Binary Code to win if $2 is bet
parameter [1:0]two_d_lose	= 2'b11;	//Binary Code to lose  if $2 is bet
//**************Parameters**************	



//**************INPUT/OUTPUT**************
	input 	clk;
	input	[5:0] seed1;
	input	[6:0] seed2;
	input	[7:0] seed3;
	output 	[3:0] rnum1, rnum2, rnum3;
	output	[1:0] bet_1d, bet_2d;
//**************INPUT/OUTPUT**************



//**************Register**************
	reg 	[1:0] bet_1d;		//register bet_1d decideds win/lose if $1 is bet 
	reg	[1:0] bet_2d;		//register bet_1d decideds win/lose if $2 is bet 
//**************Register**************



//**************Instantiation of rgen1, rgen2, and rgen3 module**************
rgen1	r1(.clk(clk), .rnum1(rnum1), .seed1(seed1));
rgen2	r2(.clk(clk), .rnum2(rnum2), .seed2(seed2));
rgen3	r3(.clk(clk), .rnum3(rnum3), .seed3(seed3));
//**************Instantiation of rgen1, rgen2, and rgen3 module**************



/*****************************Functionality******************************
***After the rnum1, rnum2, and rnum3 was created by the module rgen1, ***				
***rgen2, and rgen3, in this part they are being compared to decide   ***
***what wins or loses for $1 bet or $2 bet.			      ***
*************************************************************************/
	always @(posedge clk)
		begin
			if (rnum1 == rnum2 & rnum2 == rnum3)	//If all three numbers match $1 bet and $2 bet wins	
				begin				
				bet_1d = one_d_win;
				bet_2d = two_d_win;
				end
	
			else if (rnum1 == rnum2 | rnum1 == rnum3 | rnum2 == rnum3) //If either two numbers match $2 wins
				bet_2d = two_d_win;
			else					//else $1 and $2 loses.
			begin						
				bet_1d = one_d_lose;					
				bet_2d = two_d_lose;
			end
		end
//*****************************Functionality*****************************



endmodule
